CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 80 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
49 C:\Users\Miguel\Desktop\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
58
4 LED~
171 16 536 0 1 2
10 4
0
0 0 864 270
4 LED1
-12 -20 16 -12
2 D3
-5 -30 9 -22
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
523 0 0
2
42704.6 0
0
9 Inverter~
13 156 571 0 2 22
0 7 6
0
0 0 624 180
6 74LS04
-21 -19 21 -11
4 U16A
-8 -20 20 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 19 0
1 U
6748 0 0
2
42704.6 1
0
9 Inverter~
13 155 524 0 2 22
0 8 5
0
0 0 624 180
6 74LS04
-21 -19 21 -11
4 U11F
-8 -20 20 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 14 0
1 U
6901 0 0
2
42704.6 2
0
9 2-In AND~
219 83 540 0 3 22
0 6 5 4
0
0 0 624 180
6 74LS08
-21 -24 21 -16
4 U15D
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 18 0
1 U
842 0 0
2
42704.6 3
0
4 LED~
171 23 394 0 1 2
10 7
0
0 0 864 270
4 LED1
-12 -20 16 -12
2 D2
-5 -30 9 -22
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3277 0 0
2
42704.6 4
0
4 LED~
171 22 203 0 1 2
10 8
0
0 0 864 270
4 LED1
-12 -20 16 -12
2 D1
-5 -30 9 -22
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
4212 0 0
2
42704.6 5
0
9 2-In AND~
219 1156 136 0 3 22
0 46 21 19
0
0 0 624 180
6 74LS08
-21 -24 21 -16
4 U15C
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 18 0
1 U
4720 0 0
2
42704.6 6
0
12 SPDT Switch~
164 1293 57 0 3 11
0 46 9 46
0
0 0 4720 270
0
2 S8
9 -4 23 4
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
5551 0 0
2
42704.6 7
0
12 SPDT Switch~
164 1265 57 0 3 11
0 46 9 46
0
0 0 4720 270
0
2 S7
9 -4 23 4
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
6986 0 0
2
42704.6 8
0
9 Inverter~
13 1324 88 0 2 22
0 46 21
0
0 0 624 270
6 74LS04
-21 -19 21 -11
4 U11E
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 14 0
1 U
8745 0 0
2
42704.6 9
0
9 Inverter~
13 1214 99 0 2 22
0 46 12
0
0 0 624 270
6 74LS04
-21 -19 21 -11
4 U11D
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 14 0
1 U
9592 0 0
2
42704.6 10
0
9 2-In AND~
219 1154 190 0 3 22
0 46 46 18
0
0 0 624 180
6 74LS08
-21 -24 21 -16
4 U15B
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 18 0
1 U
8748 0 0
2
42704.6 11
0
9 2-In AND~
219 1153 240 0 3 22
0 46 21 17
0
0 0 624 180
6 74LS08
-21 -24 21 -16
4 U15A
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 18 0
1 U
7168 0 0
2
42704.6 12
0
8 3-In OR~
219 1063 190 0 4 22
0 17 18 19 11
0
0 0 624 180
4 4075
-14 -24 14 -16
4 U14B
-2 -25 26 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 17 0
1 U
631 0 0
2
42704.6 13
0
9 2-In AND~
219 1157 327 0 3 22
0 46 12 16
0
0 0 624 180
6 74LS08
-21 -24 21 -16
4 U13D
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 16 0
1 U
9466 0 0
2
42704.6 14
0
9 2-In AND~
219 1158 379 0 3 22
0 46 46 15
0
0 0 624 180
6 74LS08
-21 -24 21 -16
4 U13C
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 16 0
1 U
3266 0 0
2
42704.6 15
0
9 2-In AND~
219 1157 434 0 3 22
0 12 46 14
0
0 0 624 180
6 74LS08
-21 -24 21 -16
4 U13B
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 16 0
1 U
7693 0 0
2
42704.6 16
0
8 3-In OR~
219 1076 379 0 4 22
0 14 15 16 10
0
0 0 624 180
4 4075
-14 -24 14 -16
4 U14A
-2 -25 26 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 17 0
1 U
3723 0 0
2
42704.6 17
0
7 Ground~
168 1412 93 0 1 3
0 46
0
0 0 53360 180
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3440 0 0
2
42704.6 18
0
7 Ground~
168 1390 288 0 1 3
0 46
0
0 0 53360 180
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6263 0 0
2
42704.6 19
0
9 2-In AND~
219 178 149 0 3 22
0 23 32 31
0
0 0 624 180
6 74LS08
-21 -24 21 -16
4 U13A
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 16 0
1 U
4900 0 0
2
42704.6 20
0
12 SPDT Switch~
164 315 70 0 3 11
0 46 9 46
0
0 0 4720 270
0
2 S4
9 -4 23 4
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
8783 0 0
2
42704.6 21
0
12 SPDT Switch~
164 287 70 0 3 11
0 46 9 46
0
0 0 4720 270
0
2 S3
9 -4 23 4
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
3221 0 0
2
42704.6 22
0
9 Inverter~
13 346 101 0 2 22
0 46 32
0
0 0 624 270
6 74LS04
-21 -19 21 -11
4 U11C
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 14 0
1 U
3215 0 0
2
42704.6 23
0
9 Inverter~
13 236 112 0 2 22
0 46 24
0
0 0 624 270
6 74LS04
-21 -19 21 -11
4 U11B
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 14 0
1 U
7903 0 0
2
42704.6 24
0
9 2-In AND~
219 176 203 0 3 22
0 23 46 30
0
0 0 624 180
6 74LS08
-21 -24 21 -16
4 U12D
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 15 0
1 U
7121 0 0
2
42704.6 25
0
9 2-In AND~
219 175 253 0 3 22
0 46 32 29
0
0 0 624 180
6 74LS08
-21 -24 21 -16
4 U12C
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 15 0
1 U
4484 0 0
2
42704.6 26
0
8 3-In OR~
219 85 203 0 4 22
0 29 30 31 8
0
0 0 624 180
4 4075
-14 -24 14 -16
3 U9C
1 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 12 0
1 U
5996 0 0
2
42704.6 27
0
9 2-In AND~
219 179 340 0 3 22
0 22 24 28
0
0 0 624 180
6 74LS08
-21 -24 21 -16
4 U12B
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 15 0
1 U
7804 0 0
2
42704.6 28
0
9 2-In AND~
219 180 392 0 3 22
0 46 22 27
0
0 0 624 180
6 74LS08
-21 -24 21 -16
4 U12A
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 15 0
1 U
5523 0 0
2
42704.6 29
0
9 2-In AND~
219 179 447 0 3 22
0 24 46 26
0
0 0 624 180
6 74LS08
-21 -24 21 -16
4 U10D
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 13 0
1 U
3330 0 0
2
42704.6 30
0
8 3-In OR~
219 98 392 0 4 22
0 26 27 28 7
0
0 0 624 180
4 4075
-14 -24 14 -16
3 U9B
1 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 12 0
1 U
3465 0 0
2
42704.6 31
0
9 2-In AND~
219 481 143 0 3 22
0 34 44 42
0
0 0 624 180
6 74LS08
-21 -24 21 -16
4 U10C
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 13 0
1 U
8396 0 0
2
42704.6 32
0
12 SPDT Switch~
164 637 65 0 3 11
0 46 9 46
0
0 0 4720 270
0
2 S2
9 -4 23 4
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
3685 0 0
2
42704.6 33
0
12 SPDT Switch~
164 590 64 0 3 11
0 46 9 46
0
0 0 4720 270
0
2 S1
9 -4 23 4
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
7849 0 0
2
42704.6 34
0
9 Inverter~
13 655 97 0 2 22
0 46 44
0
0 0 624 270
6 74LS04
-21 -19 21 -11
4 U11A
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 14 0
1 U
6343 0 0
2
42704.6 35
0
9 Inverter~
13 539 106 0 2 22
0 46 35
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U7F
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 9 0
1 U
7376 0 0
2
42704.6 36
0
9 2-In AND~
219 479 197 0 3 22
0 34 46 41
0
0 0 624 180
6 74LS08
-21 -24 21 -16
4 U10B
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 13 0
1 U
9156 0 0
2
42704.6 37
0
9 2-In AND~
219 478 247 0 3 22
0 46 44 40
0
0 0 624 180
6 74LS08
-21 -24 21 -16
4 U10A
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 13 0
1 U
5776 0 0
2
42704.6 38
0
8 3-In OR~
219 388 197 0 4 22
0 40 41 42 23
0
0 0 624 180
4 4075
-14 -24 14 -16
3 U9A
1 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 12 0
1 U
7207 0 0
2
42704.6 39
0
9 2-In AND~
219 482 334 0 3 22
0 33 35 39
0
0 0 624 180
6 74LS08
-21 -24 21 -16
3 U6A
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
4459 0 0
2
42704.6 40
0
9 2-In AND~
219 483 386 0 3 22
0 46 33 38
0
0 0 624 180
6 74LS08
-21 -24 21 -16
3 U2A
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
3760 0 0
2
42704.6 41
0
9 2-In AND~
219 482 441 0 3 22
0 35 46 37
0
0 0 624 180
6 74LS08
-21 -24 21 -16
3 U1A
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
754 0 0
2
42704.6 42
0
8 3-In OR~
219 401 386 0 4 22
0 37 38 39 22
0
0 0 624 180
4 4075
-14 -24 14 -16
3 U8C
1 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 11 0
1 U
9767 0 0
2
42704.6 43
0
8 3-In OR~
219 756 393 0 4 22
0 47 48 49 33
0
0 0 624 180
4 4075
-14 -24 14 -16
3 U8B
1 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 11 0
1 U
7978 0 0
2
42704.6 44
0
9 2-In AND~
219 817 448 0 3 22
0 45 46 47
0
0 0 624 180
6 74LS08
-21 -24 21 -16
3 U5D
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 10 0
1 U
3142 0 0
2
42704.6 45
0
9 2-In AND~
219 818 393 0 3 22
0 46 10 48
0
0 0 624 180
6 74LS08
-21 -24 21 -16
3 U5C
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 10 0
1 U
3284 0 0
2
42704.6 46
0
9 2-In AND~
219 817 341 0 3 22
0 10 45 49
0
0 0 624 180
6 74LS08
-21 -24 21 -16
3 U5B
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 10 0
1 U
659 0 0
2
42704.6 47
0
8 3-In OR~
219 750 204 0 4 22
0 50 51 52 34
0
0 0 624 180
4 4075
-14 -24 14 -16
3 U8A
1 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 11 0
1 U
3800 0 0
2
42704.6 48
0
9 2-In AND~
219 813 254 0 3 22
0 46 54 50
0
0 0 624 180
6 74LS08
-21 -24 21 -16
3 U5A
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 10 0
1 U
6792 0 0
2
42704.6 49
0
9 2-In AND~
219 814 204 0 3 22
0 11 46 51
0
0 0 624 180
6 74LS08
-21 -24 21 -16
3 U3A
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
3701 0 0
2
42704.6 50
0
9 Inverter~
13 874 113 0 2 22
0 46 45
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U7E
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 9 0
1 U
6316 0 0
2
42704.6 51
0
9 Inverter~
13 984 102 0 2 22
0 46 54
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U7A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 9 0
1 U
8734 0 0
2
5.89779e-315 0
0
12 SPDT Switch~
164 925 71 0 3 11
0 46 9 46
0
0 0 4720 270
0
2 S6
9 -4 23 4
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
7988 0 0
2
42704.6 52
0
12 SPDT Switch~
164 953 71 0 3 11
0 46 9 46
0
0 0 4720 270
0
2 S5
9 -4 23 4
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
3217 0 0
2
42704.6 53
0
9 2-In AND~
219 816 150 0 3 22
0 11 54 52
0
0 0 624 180
6 74LS08
-21 -24 21 -16
3 U4B
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
3965 0 0
2
42704.6 54
0
7 Ground~
168 43 102 0 1 3
0 46
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8239 0 0
2
42704.6 55
0
2 +V
167 42 39 0 1 3
0 9
0
0 0 54256 0
3 10V
-11 -24 10 -16
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
828 0 0
2
42704.6 56
0
119
2 0 46 0 0 4096 3 26 0 0 64 2
194 194
286 194
2 0 46 0 0 4096 2 16 0 0 3 3
1176 370
1390 370
1390 336
1 1 46 0 0 4096 2 15 20 0 0 3
1175 336
1390 336
1390 296
1 0 46 0 0 4096 2 12 0 0 5 3
1172 199
1412 199
1412 145
1 1 46 0 0 0 2 7 19 0 0 3
1174 145
1412 145
1412 101
3 1 4 0 0 4224 0 4 1 0 0 4
56 540
36 540
36 534
28 534
2 2 5 0 0 4224 0 3 4 0 0 4
140 524
111 524
111 531
101 531
2 1 6 0 0 4224 0 2 4 0 0 4
141 571
111 571
111 549
101 549
0 1 7 0 0 8320 0 0 2 15 0 5
63 392
63 504
190 504
190 571
177 571
0 1 8 0 0 4224 0 0 3 16 0 5
44 201
44 509
184 509
184 524
176 524
2 0 9 0 0 4096 0 22 0 0 117 2
318 54
318 34
3 0 46 0 0 0 2 22 0 0 119 2
310 54
310 39
2 0 9 0 0 0 0 23 0 0 117 2
290 54
290 34
3 0 46 0 0 0 2 23 0 0 119 2
282 54
282 39
1 4 7 0 0 0 0 5 32 0 0 4
35 392
77 392
77 392
71 392
1 4 8 0 0 0 0 6 28 0 0 4
34 201
64 201
64 203
58 203
0 3 46 0 0 0 2 0 9 18 0 2
1260 22
1260 41
0 3 46 0 0 8192 2 0 8 119 0 4
945 39
945 22
1288 22
1288 41
0 2 9 0 0 0 0 0 9 20 0 2
1268 27
1268 41
0 2 9 0 0 8192 0 0 8 117 0 4
956 34
956 27
1296 27
1296 41
2 4 10 0 0 4096 0 47 18 0 0 4
836 384
1050 384
1050 379
1049 379
1 4 10 0 0 4224 0 48 18 0 0 4
835 350
1055 350
1055 379
1049 379
1 4 11 0 0 4096 0 51 14 0 0 4
832 213
1037 213
1037 190
1036 190
1 4 11 0 0 4224 0 56 14 0 0 4
834 159
1042 159
1042 190
1036 190
0 1 12 0 0 4096 0 0 17 39 0 4
1217 444
1185 444
1185 443
1175 443
0 2 46 0 0 4096 13 0 17 43 0 2
1292 425
1175 425
0 1 46 0 0 0 13 0 16 43 0 2
1292 388
1176 388
2 0 12 0 0 4096 0 15 0 0 39 2
1175 318
1217 318
1 3 14 0 0 8320 0 18 17 0 0 4
1095 388
1124 388
1124 434
1130 434
2 3 15 0 0 4224 0 18 16 0 0 2
1094 379
1131 379
3 3 16 0 0 8320 0 18 15 0 0 4
1095 370
1124 370
1124 327
1130 327
1 3 17 0 0 8320 0 14 13 0 0 4
1082 199
1120 199
1120 240
1126 240
2 3 18 0 0 4224 0 14 12 0 0 2
1081 190
1127 190
3 3 19 0 0 8320 0 14 7 0 0 4
1082 181
1123 181
1123 136
1129 136
0 1 46 0 0 4096 20 0 13 41 0 2
1264 249
1171 249
0 2 21 0 0 4096 0 0 13 42 0 2
1327 231
1171 231
2 0 46 0 0 0 20 12 0 0 41 2
1172 181
1264 181
0 2 21 0 0 0 0 0 7 42 0 2
1327 127
1174 127
2 0 12 0 0 4224 0 11 0 0 0 2
1217 117
1217 521
1 1 46 0 0 0 20 9 11 0 0 4
1264 75
1264 78
1217 78
1217 81
1 0 46 0 0 4224 20 9 0 0 0 2
1264 75
1264 522
2 0 21 0 0 4224 0 10 0 0 0 2
1327 106
1327 522
1 0 46 0 0 4224 13 8 0 0 0 2
1292 75
1292 522
1 1 46 0 0 0 13 8 10 0 0 3
1292 75
1292 70
1327 70
2 4 22 0 0 4096 0 30 44 0 0 4
198 383
375 383
375 386
374 386
1 4 22 0 0 4224 0 29 44 0 0 4
197 349
380 349
380 386
374 386
1 4 23 0 0 4096 0 26 40 0 0 4
194 212
362 212
362 197
361 197
1 4 23 0 0 4224 0 21 40 0 0 4
196 158
367 158
367 197
361 197
0 1 24 0 0 4096 0 0 31 62 0 2
239 456
197 456
0 2 46 0 0 4096 25 0 31 66 0 2
314 438
197 438
0 1 46 0 0 0 25 0 30 66 0 2
314 401
198 401
2 0 24 0 0 0 0 29 0 0 62 2
197 331
239 331
1 3 26 0 0 8320 0 32 31 0 0 4
117 401
146 401
146 447
152 447
2 3 27 0 0 4224 0 32 30 0 0 2
116 392
153 392
3 3 28 0 0 8320 0 32 29 0 0 4
117 383
146 383
146 340
152 340
1 3 29 0 0 8320 0 28 27 0 0 4
104 212
142 212
142 253
148 253
2 3 30 0 0 4224 0 28 26 0 0 2
103 203
149 203
3 3 31 0 0 8320 0 28 21 0 0 4
104 194
145 194
145 149
151 149
0 1 46 0 0 4096 3 0 27 64 0 2
286 262
193 262
0 2 32 0 0 4096 0 0 27 65 0 2
349 244
193 244
0 2 32 0 0 0 0 0 21 65 0 2
349 140
196 140
2 0 24 0 0 4224 0 25 0 0 0 2
239 130
239 534
1 1 46 0 0 0 3 23 25 0 0 4
286 88
286 91
239 91
239 94
1 0 46 0 0 4224 3 23 0 0 0 2
286 88
286 535
2 0 32 0 0 4224 0 24 0 0 0 2
349 119
349 535
1 0 46 0 0 4224 25 22 0 0 0 2
314 88
314 535
1 1 46 0 0 0 25 22 24 0 0 3
314 88
314 83
349 83
0 3 46 0 0 0 2 0 35 119 0 3
582 39
582 48
585 48
0 2 9 0 0 0 0 0 35 117 0 2
593 34
593 48
0 3 46 0 0 0 2 0 34 119 0 3
611 39
611 49
632 49
0 2 9 0 0 0 0 0 34 117 0 4
621 34
621 41
640 41
640 49
2 4 33 0 0 4096 0 42 45 0 0 4
501 377
710 377
710 393
729 393
1 4 33 0 0 4224 0 41 45 0 0 4
500 343
715 343
715 393
729 393
1 4 34 0 0 4096 0 38 49 0 0 4
497 206
697 206
697 204
723 204
1 4 34 0 0 4224 0 33 49 0 0 4
499 152
702 152
702 204
723 204
0 1 35 0 0 4096 0 0 43 90 0 2
542 450
500 450
0 2 46 0 0 4096 36 0 43 94 0 2
617 432
500 432
0 1 46 0 0 0 36 0 42 94 0 2
617 395
501 395
2 0 35 0 0 0 0 41 0 0 90 2
500 325
542 325
1 3 37 0 0 8320 0 44 43 0 0 4
420 395
449 395
449 441
455 441
2 3 38 0 0 4224 0 44 42 0 0 2
419 386
456 386
3 3 39 0 0 8320 0 44 41 0 0 4
420 377
449 377
449 334
455 334
1 3 40 0 0 8320 0 40 39 0 0 4
407 206
445 206
445 247
451 247
2 3 41 0 0 4224 0 40 38 0 0 2
406 197
452 197
3 3 42 0 0 8320 0 40 33 0 0 4
407 188
448 188
448 143
454 143
0 1 46 0 0 4096 43 0 39 92 0 2
589 256
496 256
0 2 44 0 0 4096 0 0 39 93 0 2
652 238
496 238
2 0 46 0 0 0 43 38 0 0 92 2
497 188
589 188
0 2 44 0 0 0 0 0 33 93 0 2
652 134
499 134
2 0 35 0 0 4224 0 37 0 0 0 2
542 124
542 528
1 1 46 0 0 0 43 35 37 0 0 4
589 82
589 85
542 85
542 88
1 0 46 0 0 4224 43 35 0 0 0 2
589 82
589 529
2 0 44 0 0 12416 0 36 0 0 0 4
658 115
658 134
652 134
652 529
1 0 46 0 0 4224 36 34 0 0 0 4
636 83
636 395
617 395
617 529
1 1 46 0 0 0 36 34 36 0 0 3
636 83
636 79
658 79
0 1 45 0 0 4096 0 0 46 110 0 2
877 457
835 457
0 2 46 0 0 4096 0 0 46 114 0 2
952 439
835 439
0 1 46 0 0 0 0 0 47 114 0 2
952 402
836 402
2 0 45 0 0 0 0 48 0 0 110 2
835 332
877 332
1 3 47 0 0 8320 0 45 46 0 0 4
775 402
784 402
784 448
790 448
2 3 48 0 0 4224 0 45 47 0 0 2
774 393
791 393
3 3 49 0 0 8320 0 45 48 0 0 4
775 384
784 384
784 341
790 341
1 3 50 0 0 8320 0 49 50 0 0 4
769 213
780 213
780 254
786 254
2 3 51 0 0 4224 0 49 51 0 0 2
768 204
787 204
3 3 52 0 0 8320 0 49 56 0 0 4
769 195
783 195
783 150
789 150
0 1 46 0 0 4096 53 0 50 112 0 2
924 263
831 263
0 2 54 0 0 4096 0 0 50 113 0 2
987 245
831 245
2 0 46 0 0 0 53 51 0 0 112 2
832 195
924 195
0 2 54 0 0 0 0 0 56 113 0 2
987 141
834 141
2 0 45 0 0 4224 0 52 0 0 0 2
877 131
877 535
1 1 46 0 0 0 53 54 52 0 0 4
924 89
924 92
877 92
877 95
1 0 46 0 0 4224 53 54 0 0 0 2
924 89
924 536
2 0 54 0 0 4224 0 53 0 0 0 2
987 120
987 536
1 0 46 0 0 4224 0 55 0 0 0 2
952 89
952 536
1 1 46 0 0 0 0 55 53 0 0 3
952 89
952 84
987 84
0 2 9 0 0 0 0 0 54 117 0 2
928 34
928 55
1 2 9 0 0 16512 0 58 55 0 0 6
42 48
42 57
214 57
214 34
956 34
956 55
0 3 46 0 0 0 2 0 54 119 0 2
920 39
920 55
1 3 46 0 0 16512 2 57 55 0 0 6
43 96
43 71
219 71
219 39
948 39
948 55
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
