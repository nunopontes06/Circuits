CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1918 1059
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
5 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
44
6 74136~
219 244 195 0 3 22
0 5 35 8
0
0 0 608 270
7 74LS136
-24 -24 25 -16
3 U6A
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
5130 0 0
2
44200.9 0
0
6 74136~
219 421 189 0 3 22
0 5 6 9
0
0 0 608 270
7 74LS136
-24 -24 25 -16
3 U7D
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 7 0
1 U
391 0 0
2
44200.9 1
0
6 74136~
219 580 186 0 3 22
0 5 36 10
0
0 0 608 270
7 74LS136
-24 -24 25 -16
3 U7C
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 7 0
1 U
3124 0 0
2
44200.9 2
0
6 74136~
219 967 201 0 3 22
0 2 5 3
0
0 0 608 180
7 74LS136
-24 -24 25 -16
3 U7B
-2 -25 19 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
3421 0 0
2
44200.9 3
0
2 +V
167 1090 111 0 1 3
0 7
0
0 0 54240 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8157 0 0
2
44200.9 4
0
7 Ground~
168 1047 266 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5572 0 0
2
44200.9 5
0
12 SPDT Switch~
164 1019 194 0 3 11
0 5 2 7
0
0 0 4704 180
0
2 S9
-7 -16 7 -8
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
8901 0 0
2
44200.9 6
0
6 74136~
219 765 237 0 3 22
0 5 37 11
0
0 0 608 270
7 74LS136
-24 -24 25 -16
3 U7A
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
7361 0 0
2
44200.9 7
0
6 74136~
219 818 416 0 3 22
0 12 11 32
0
0 0 608 270
7 74LS136
-24 -24 25 -16
3 U1A
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
4747 0 0
2
44200.9 8
0
9 2-In AND~
219 760 418 0 3 22
0 11 12 34
0
0 0 608 270
6 74LS08
-21 -24 21 -16
3 U2A
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
972 0 0
2
44200.9 9
0
9 2-In AND~
219 772 548 0 3 22
0 3 32 33
0
0 0 608 270
6 74LS08
-21 -24 21 -16
3 U2B
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
3472 0 0
2
44200.9 10
0
6 74136~
219 827 556 0 3 22
0 3 32 31
0
0 0 608 270
7 74LS136
-24 -24 25 -16
3 U1B
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
9998 0 0
2
44200.9 11
0
8 2-In OR~
219 746 676 0 3 22
0 33 34 15
0
0 0 608 270
6 74LS32
-21 -24 21 -16
3 U3A
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3536 0 0
2
44200.9 12
0
4 LED~
171 830 927 0 2 2
10 31 2
0
0 0 864 0
4 LED1
17 0 45 8
2 D1
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
4597 0 0
2
44200.9 13
0
4 LED~
171 653 935 0 2 2
10 26 2
0
0 0 864 0
4 LED1
17 0 45 8
2 D2
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3835 0 0
2
44200.9 14
0
8 2-In OR~
219 569 684 0 3 22
0 28 29 14
0
0 0 608 270
6 74LS32
-21 -24 21 -16
3 U3B
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
3670 0 0
2
44200.9 15
0
6 74136~
219 650 564 0 3 22
0 15 27 26
0
0 0 608 270
7 74LS136
-24 -24 25 -16
3 U1C
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
5616 0 0
2
44200.9 16
0
9 2-In AND~
219 595 556 0 3 22
0 15 27 28
0
0 0 608 270
6 74LS08
-21 -24 21 -16
3 U2C
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
9323 0 0
2
44200.9 17
0
9 2-In AND~
219 583 426 0 3 22
0 10 30 29
0
0 0 608 270
6 74LS08
-21 -24 21 -16
3 U2D
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
317 0 0
2
44200.9 18
0
6 74136~
219 641 424 0 3 22
0 10 30 27
0
0 0 608 270
7 74LS136
-24 -24 25 -16
3 U1D
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
3108 0 0
2
44200.9 19
0
4 LED~
171 489 931 0 2 2
10 21 2
0
0 0 864 0
4 LED1
17 0 45 8
2 D3
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
4299 0 0
2
44200.9 20
0
8 2-In OR~
219 405 680 0 3 22
0 23 24 13
0
0 0 608 270
6 74LS32
-21 -24 21 -16
3 U3C
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
9672 0 0
2
44200.9 21
0
6 74136~
219 486 560 0 3 22
0 14 22 21
0
0 0 608 270
7 74LS136
-24 -24 25 -16
3 U4A
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
7876 0 0
2
44200.9 22
0
9 2-In AND~
219 431 552 0 3 22
0 14 22 23
0
0 0 608 270
6 74LS08
-21 -24 21 -16
3 U5A
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
6369 0 0
2
44200.9 23
0
9 2-In AND~
219 419 422 0 3 22
0 9 25 24
0
0 0 608 270
6 74LS08
-21 -24 21 -16
3 U5B
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
9172 0 0
2
44200.9 24
0
6 74136~
219 477 420 0 3 22
0 9 25 22
0
0 0 608 270
7 74LS136
-24 -24 25 -16
3 U4B
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
7100 0 0
2
44200.9 25
0
4 LED~
171 313 941 0 2 2
10 17 2
0
0 0 864 0
4 LED1
17 0 45 8
2 D4
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3820 0 0
2
44200.9 26
0
8 2-In OR~
219 229 690 0 3 22
0 19 20 16
0
0 0 608 270
6 74LS32
-21 -24 21 -16
3 U3D
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
7678 0 0
2
44200.9 27
0
6 74136~
219 310 570 0 3 22
0 13 18 17
0
0 0 608 270
7 74LS136
-24 -24 25 -16
3 U4C
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
961 0 0
2
44200.9 28
0
9 2-In AND~
219 255 562 0 3 22
0 13 18 19
0
0 0 608 270
6 74LS08
-21 -24 21 -16
3 U5C
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
3178 0 0
2
44200.9 29
0
9 2-In AND~
219 243 432 0 3 22
0 8 4 20
0
0 0 608 270
6 74LS08
-21 -24 21 -16
3 U5D
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
3409 0 0
2
44200.9 30
0
6 74136~
219 301 430 0 3 22
0 8 4 18
0
0 0 608 270
7 74LS136
-24 -24 25 -16
3 U4D
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
3951 0 0
2
44200.9 31
0
4 LED~
171 232 936 0 2 2
10 16 2
0
0 0 864 0
4 LED1
17 0 45 8
2 D5
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
8885 0 0
2
44200.9 32
0
7 Ground~
168 466 1045 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3780 0 0
2
44200.9 33
0
12 SPDT Switch~
164 219 93 0 10 11
0 4 2 38 0 0 0 0 0 0
1
0
0 0 4704 270
0
2 S8
1 17 15 25
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
9265 0 0
2
5.89699e-315 0
0
12 SPDT Switch~
164 238 96 0 10 11
0 35 2 38 0 0 0 0 0 0
1
0
0 0 4704 270
0
2 S7
5 15 19 23
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
9442 0 0
2
5.89699e-315 5.26354e-315
0
12 SPDT Switch~
164 395 83 0 10 11
0 25 2 38 0 0 0 0 0 0
1
0
0 0 4704 270
0
2 S6
1 17 15 25
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
9424 0 0
2
5.89699e-315 5.30499e-315
0
12 SPDT Switch~
164 414 86 0 10 11
0 6 2 38 0 0 0 0 0 0
1
0
0 0 4704 270
0
2 S5
5 15 19 23
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
9968 0 0
2
5.89699e-315 5.32571e-315
0
12 SPDT Switch~
164 559 87 0 10 11
0 30 2 38 0 0 0 0 0 0
1
0
0 0 4704 270
0
2 S4
1 17 15 25
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
9281 0 0
2
5.89699e-315 5.34643e-315
0
12 SPDT Switch~
164 578 90 0 10 11
0 36 2 38 0 0 0 0 0 0
1
0
0 0 4704 270
0
2 S3
5 15 19 23
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
8464 0 0
2
5.89699e-315 5.3568e-315
0
12 SPDT Switch~
164 755 82 0 10 11
0 37 2 38 0 0 0 0 0 0
1
0
0 0 4704 270
0
2 S2
5 15 19 23
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
7168 0 0
2
5.89699e-315 5.36716e-315
0
12 SPDT Switch~
164 736 79 0 10 11
0 12 2 38 0 0 0 0 0 0
1
0
0 0 4704 270
0
2 S1
1 17 15 25
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
3171 0 0
2
5.89699e-315 5.37752e-315
0
2 +V
167 962 33 0 1 3
0 38
0
0 0 54240 0
3 10V
-11 -22 10 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4139 0 0
2
5.89699e-315 5.38788e-315
0
7 Ground~
168 65 81 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6435 0 0
2
44200.9 34
0
79
1 0 3 0 0 8192 0 11 0 0 2 3
779 526
779 515
839 515
1 3 3 0 0 12416 0 12 4 0 0 5
839 537
839 445
942 445
942 201
940 201
0 2 4 0 0 4096 0 0 32 4 0 3
218 361
295 361
295 411
1 2 4 0 0 4224 0 35 31 0 0 4
218 111
218 409
232 409
232 410
1 0 5 0 0 4096 0 8 0 0 8 2
777 218
777 142
1 0 5 0 0 0 0 3 0 0 8 2
592 167
592 142
1 0 5 0 0 0 0 2 0 0 8 2
433 170
433 142
1 1 5 0 0 8320 0 7 1 0 0 4
1002 192
1002 142
256 142
256 176
0 2 6 0 0 8320 0 0 2 61 0 3
413 107
415 107
415 170
1 0 2 0 0 4096 0 4 0 0 12 2
989 210
1047 210
2 1 5 0 0 0 0 4 7 0 0 2
989 192
1002 192
1 2 2 0 0 4096 0 6 7 0 0 3
1047 260
1047 196
1036 196
1 3 7 0 0 4224 0 5 7 0 0 3
1090 120
1090 188
1036 188
0 1 8 0 0 4096 0 0 32 15 0 3
250 396
313 396
313 411
3 1 8 0 0 4224 0 1 31 0 0 4
247 225
247 382
250 382
250 410
0 1 9 0 0 4096 0 0 26 17 0 3
426 387
489 387
489 401
3 1 9 0 0 4224 0 2 25 0 0 4
424 219
424 370
426 370
426 400
0 1 10 0 0 4096 0 0 20 19 0 3
590 395
653 395
653 405
3 1 10 0 0 4224 0 3 19 0 0 4
583 216
583 375
590 375
590 404
0 2 11 0 0 4096 0 0 9 22 0 3
767 388
812 388
812 397
0 1 12 0 0 4096 0 0 9 59 0 3
735 372
830 372
830 397
3 1 11 0 0 4224 0 8 10 0 0 4
768 267
768 375
767 375
767 396
1 0 13 0 0 8192 0 30 0 0 32 3
262 540
262 531
322 531
1 0 14 0 0 8192 0 24 0 0 33 3
438 530
438 522
498 522
1 0 15 0 0 8192 0 18 0 0 34 3
602 534
602 527
662 527
0 1 2 0 0 0 2 0 34 30 0 2
466 1002
466 1039
2 0 2 0 0 0 2 15 0 0 30 2
653 945
653 1002
2 0 2 0 0 0 2 21 0 0 30 2
489 941
489 1002
2 0 2 0 0 0 2 27 0 0 30 2
313 951
313 1002
2 2 2 0 0 8192 2 14 33 0 0 4
830 937
830 1002
232 1002
232 946
3 1 16 0 0 4224 0 28 33 0 0 2
232 720
232 926
3 1 13 0 0 12416 0 22 29 0 0 6
408 710
408 727
368 727
368 504
322 504
322 551
1 3 14 0 0 12416 0 23 16 0 0 6
498 541
498 499
539 499
539 728
572 728
572 714
3 1 15 0 0 12416 0 13 17 0 0 6
749 706
749 730
707 730
707 501
662 501
662 545
3 1 17 0 0 4224 0 29 27 0 0 2
313 600
313 931
2 0 18 0 0 4096 0 30 0 0 37 3
244 540
244 480
304 480
3 2 18 0 0 4224 0 32 29 0 0 2
304 460
304 551
3 1 19 0 0 4224 0 30 28 0 0 4
253 585
253 659
241 659
241 674
3 2 20 0 0 8320 0 31 28 0 0 3
241 455
223 455
223 674
3 1 21 0 0 4224 0 23 21 0 0 2
489 590
489 921
2 0 22 0 0 4096 0 24 0 0 42 3
420 530
420 470
480 470
3 2 22 0 0 4224 0 26 23 0 0 2
480 450
480 541
3 1 23 0 0 4224 0 24 22 0 0 4
429 575
429 649
417 649
417 664
3 2 24 0 0 8320 0 25 22 0 0 3
417 445
399 445
399 664
2 0 25 0 0 8192 26 26 0 0 46 3
471 401
471 379
394 379
1 2 25 0 0 4224 26 37 25 0 0 3
394 101
394 400
408 400
3 1 26 0 0 4224 0 17 15 0 0 2
653 594
653 925
2 0 27 0 0 4096 0 18 0 0 49 3
584 534
584 474
644 474
3 2 27 0 0 4224 0 20 17 0 0 2
644 454
644 545
3 1 28 0 0 4224 0 18 16 0 0 4
593 579
593 653
581 653
581 668
3 2 29 0 0 8320 0 19 16 0 0 3
581 449
563 449
563 668
2 0 30 0 0 8192 31 20 0 0 53 3
635 405
635 383
558 383
1 2 30 0 0 4224 31 39 19 0 0 3
558 105
558 404
572 404
3 1 31 0 0 4224 0 12 14 0 0 2
830 586
830 917
2 0 32 0 0 4096 0 11 0 0 56 3
761 526
761 466
821 466
3 2 32 0 0 4224 0 9 12 0 0 2
821 446
821 537
3 1 33 0 0 4224 0 11 13 0 0 4
770 571
770 645
758 645
758 660
3 2 34 0 0 8320 0 10 13 0 0 3
758 441
740 441
740 660
1 2 12 0 0 4224 0 42 10 0 0 3
735 97
735 396
749 396
1 2 35 0 0 12416 5 36 1 0 0 4
237 114
237 124
238 124
238 176
1 0 6 0 0 0 7 38 0 0 0 2
413 104
413 112
1 2 36 0 0 12416 9 40 3 0 0 4
577 108
577 117
574 117
574 167
1 2 37 0 0 12416 12 41 8 0 0 4
754 100
754 112
759 112
759 218
2 0 2 0 0 0 2 42 0 0 71 2
739 63
739 34
2 0 2 0 0 0 2 40 0 0 71 2
581 74
581 34
2 0 2 0 0 0 2 39 0 0 71 2
562 71
562 34
2 0 2 0 0 0 2 38 0 0 71 2
417 70
417 34
2 0 2 0 0 0 2 37 0 0 71 2
398 67
398 34
2 0 2 0 0 0 2 36 0 0 71 2
241 80
241 34
2 0 2 0 0 0 2 35 0 0 71 2
222 77
222 34
1 2 2 0 0 8320 2 44 41 0 0 4
65 75
65 34
758 34
758 66
3 0 38 0 0 4096 3 36 0 0 79 2
233 80
233 45
3 0 38 0 0 0 3 38 0 0 79 2
409 70
409 45
3 0 38 0 0 0 3 41 0 0 79 2
750 66
750 45
3 0 38 0 0 0 3 40 0 0 79 2
573 74
573 45
3 0 38 0 0 0 3 42 0 0 79 2
731 63
731 45
3 0 38 0 0 0 3 39 0 0 79 2
554 71
554 45
3 0 38 0 0 0 3 37 0 0 79 2
390 67
390 45
1 3 38 0 0 8320 3 43 35 0 0 4
962 42
962 45
214 45
214 77
8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
398 4 437 28
409 13 425 29
2 A2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
731 5 770 29
742 14 758 30
2 A0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
711 5 750 29
722 14 738 30
2 B0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
560 6 599 30
571 15 587 31
2 A1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
540 5 579 29
551 14 567 30
2 B1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
376 4 415 28
387 13 403 29
2 B2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
201 4 240 28
212 13 228 29
2 B3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
225 4 264 28
236 13 252 29
2 A3
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
