CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
58 C:\Users\joaop\Desktop\circuitmaker+traxmaker+2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
45
7 Ground~
168 1165 352 0 1 3
0 0
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5130 0 0
2
43084.4 0
0
9 Inverter~
13 994 333 0 2 22
0 4 3
0
0 0 608 180
6 74LS04
-21 -19 21 -11
3 U7B
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 8 0
1 U
391 0 0
2
43084.4 0
0
9 Inverter~
13 704 331 0 2 22
0 6 5
0
0 0 608 180
6 74LS04
-21 -19 21 -11
3 U7A
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 8 0
1 U
3124 0 0
2
43084.4 1
0
9 Inverter~
13 434 320 0 2 22
0 8 7
0
0 0 608 180
6 74LS04
-21 -19 21 -11
3 U1F
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 7 0
1 U
3421 0 0
2
43084.4 2
0
9 Inverter~
13 184 322 0 2 22
0 10 9
0
0 0 608 180
6 74LS04
-21 -19 21 -11
3 U1E
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 7 0
1 U
8157 0 0
2
43084.4 3
0
9 Inverter~
13 959 230 0 2 22
0 12 11
0
0 0 608 180
6 74LS04
-21 -19 21 -11
3 U1D
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 7 0
1 U
5572 0 0
2
43084.4 4
0
9 Inverter~
13 668 215 0 2 22
0 14 13
0
0 0 608 180
6 74LS04
-21 -19 21 -11
3 U1C
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 7 0
1 U
8901 0 0
2
43084.4 5
0
9 Inverter~
13 387 220 0 2 22
0 16 15
0
0 0 608 512
6 74LS04
-21 -19 21 -11
3 U1B
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 7 0
1 U
7361 0 0
2
43084.4 6
0
9 Inverter~
13 141 217 0 2 22
0 18 17
0
0 0 608 180
6 74LS04
-21 -19 21 -11
3 U1A
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 7 0
1 U
4747 0 0
2
43084.4 7
0
4 LED~
171 43 475 0 2 2
10 20 2
0
0 0 880 0
4 LED0
17 0 45 8
2 D5
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
972 0 0
2
43084.4 8
0
7 Ground~
168 629 579 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3472 0 0
2
43084.4 9
0
4 LED~
171 258 480 0 2 2
10 24 2
0
0 0 880 0
4 LED0
17 0 45 8
2 D4
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
9998 0 0
2
43084.4 10
0
4 LED~
171 508 468 0 2 2
10 23 2
0
0 0 880 0
4 LED0
17 0 45 8
2 D3
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3536 0 0
2
43084.4 11
0
4 LED~
171 788 473 0 2 2
10 22 2
0
0 0 880 0
4 LED0
17 0 45 8
2 D2
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
4597 0 0
2
43084.4 12
0
4 LED~
171 1076 494 0 2 2
10 21 2
0
0 0 880 0
4 LED0
17 0 45 8
2 D1
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3835 0 0
2
43084.4 13
0
7 Ground~
168 78 132 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3670 0 0
2
43084.4 14
0
2 +V
167 120 62 0 1 3
0 25
0
0 0 54240 0
3 10V
-11 -23 10 -15
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5616 0 0
2
43084.4 15
0
12 SPDT Switch~
164 1090 160 0 10 11
0 31 25 2 0 0 0 0 0 0
1
0
0 0 4704 270
0
2 S8
9 -4 23 4
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
9323 0 0
2
43084.4 16
0
12 SPDT Switch~
164 999 161 0 10 11
0 12 25 2 0 0 0 0 0 0
1
0
0 0 4704 270
0
2 S7
9 -4 23 4
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
317 0 0
2
43084.4 17
0
12 SPDT Switch~
164 796 162 0 10 11
0 40 25 2 0 0 0 0 0 0
1
0
0 0 4704 270
0
2 S6
9 -4 23 4
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
3108 0 0
2
43084.4 18
0
12 SPDT Switch~
164 713 161 0 10 11
0 14 25 2 0 0 0 0 0 0
1
0
0 0 4704 270
0
2 S5
9 -4 23 4
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
4299 0 0
2
43084.4 19
0
12 SPDT Switch~
164 524 158 0 10 11
0 37 25 2 0 0 0 0 0 0
1
0
0 0 4704 270
0
2 S4
9 -4 23 4
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
9672 0 0
2
43084.4 20
0
12 SPDT Switch~
164 426 158 0 10 11
0 16 25 2 0 0 0 0 0 0
1
0
0 0 4704 270
0
2 S3
9 -4 23 4
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
7876 0 0
2
43084.4 21
0
12 SPDT Switch~
164 274 162 0 10 11
0 34 25 2 0 0 0 0 0 0
1
0
0 0 4704 270
0
2 S2
9 -4 23 4
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
6369 0 0
2
43084.4 22
0
12 SPDT Switch~
164 184 159 0 10 11
0 18 25 2 0 0 0 0 0 0
1
0
0 0 4704 270
0
2 S1
9 -4 23 4
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
9172 0 0
2
43084.4 23
0
6 74136~
219 1070 282 0 3 22
0 31 12 4
0
0 0 608 270
7 74LS136
-24 -24 25 -16
3 U6D
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 6 0
1 U
7100 0 0
2
43084.4 24
0
6 74136~
219 1071 374 0 3 22
0 19 4 21
0
0 0 608 270
7 74LS136
-24 -24 25 -16
3 U6C
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
3820 0 0
2
43084.4 25
0
9 2-In AND~
219 961 295 0 3 22
0 31 11 30
0
0 0 608 180
6 74LS08
-21 -24 21 -16
3 U5D
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
7678 0 0
2
43084.4 26
0
9 2-In AND~
219 965 418 0 3 22
0 19 3 29
0
0 0 608 180
6 74LS08
-21 -24 21 -16
3 U5C
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
961 0 0
2
43084.4 27
0
8 2-In OR~
219 889 337 0 3 22
0 29 30 28
0
0 0 608 180
6 74LS32
-21 -24 21 -16
3 U4D
1 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
3178 0 0
2
43084.4 28
0
6 74136~
219 241 272 0 3 22
0 34 18 10
0
0 0 608 270
7 74LS136
-24 -24 25 -16
3 U6B
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
3409 0 0
2
43084.4 29
0
6 74136~
219 255 360 0 3 22
0 26 10 24
0
0 0 608 270
7 74LS136
-24 -24 25 -16
3 U6A
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
3951 0 0
2
43084.4 30
0
9 2-In AND~
219 138 274 0 3 22
0 34 17 33
0
0 0 608 180
6 74LS08
-21 -24 21 -16
3 U5B
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
8885 0 0
2
43084.4 31
0
9 2-In AND~
219 164 411 0 3 22
0 26 9 32
0
0 0 608 180
6 74LS08
-21 -24 21 -16
3 U5A
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
3780 0 0
2
43084.4 32
0
8 2-In OR~
219 73 323 0 3 22
0 32 33 20
0
0 0 608 180
6 74LS32
-21 -24 21 -16
3 U4C
1 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
9265 0 0
2
43084.4 33
0
6 74136~
219 491 274 0 3 22
0 37 16 8
0
0 0 608 270
7 74LS136
-24 -24 25 -16
3 U2D
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
9442 0 0
2
43084.4 34
0
6 74136~
219 505 362 0 3 22
0 27 8 23
0
0 0 608 270
7 74LS136
-24 -24 25 -16
3 U2C
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
9424 0 0
2
43084.4 35
0
9 2-In AND~
219 396 284 0 3 22
0 37 15 36
0
0 0 608 180
6 74LS08
-21 -24 21 -16
3 U3D
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
9968 0 0
2
43084.4 36
0
9 2-In AND~
219 403 402 0 3 22
0 27 7 35
0
0 0 608 180
6 74LS08
-21 -24 21 -16
3 U3C
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
9281 0 0
2
43084.4 37
0
8 2-In OR~
219 323 325 0 3 22
0 35 36 26
0
0 0 608 180
6 74LS32
-21 -24 21 -16
3 U4B
1 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
8464 0 0
2
43084.4 38
0
8 2-In OR~
219 603 329 0 3 22
0 38 39 27
0
0 0 608 180
6 74LS32
-21 -24 21 -16
3 U4A
1 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
7168 0 0
2
43084.4 39
0
9 2-In AND~
219 689 405 0 3 22
0 28 5 38
0
0 0 608 180
6 74LS08
-21 -24 21 -16
3 U3B
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
3171 0 0
2
43084.4 40
0
9 2-In AND~
219 669 285 0 3 22
0 40 13 39
0
0 0 608 180
6 74LS08
-21 -24 21 -16
3 U3A
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
4139 0 0
2
43084.4 41
0
6 74136~
219 785 366 0 3 22
0 28 6 22
0
0 0 608 270
7 74LS136
-24 -24 25 -16
3 U2B
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
6435 0 0
2
43084.4 42
0
6 74136~
219 771 278 0 3 22
0 40 14 6
0
0 0 608 270
7 74LS136
-24 -24 25 -16
3 U2A
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
5283 0 0
2
43084.4 43
0
74
2 0 2 0 0 8192 0 14 0 0 2 5
788 483
794 483
794 500
795 500
795 504
2 0 2 0 0 4096 0 15 0 0 31 3
1076 504
628 504
628 515
2 2 3 0 0 16512 0 2 29 0 0 6
979 333
975 333
975 361
1002 361
1002 409
983 409
1 0 4 0 0 8320 0 2 0 0 14 3
1015 333
1015 320
1065 320
2 2 5 0 0 12416 0 3 42 0 0 5
689 331
689 351
719 351
719 396
707 396
1 0 6 0 0 4224 0 3 0 0 11 2
725 331
779 331
2 2 7 0 0 16512 0 4 39 0 0 6
419 320
415 320
415 352
436 352
436 393
421 393
1 0 8 0 0 4224 0 4 0 0 12 2
455 320
494 320
2 2 9 0 0 16512 0 5 34 0 0 6
169 322
162 322
162 350
186 350
186 402
182 402
0 1 10 0 0 4224 0 0 5 13 0 2
244 322
205 322
3 2 6 0 0 0 0 45 44 0 0 3
774 308
779 308
779 347
3 2 8 0 0 0 0 36 37 0 0 4
494 304
494 330
499 330
499 343
3 2 10 0 0 0 0 31 32 0 0 4
244 302
244 328
249 328
249 341
3 2 4 0 0 0 0 26 27 0 0 4
1073 312
1073 320
1065 320
1065 355
2 2 11 0 0 12416 0 6 28 0 0 6
944 230
927 230
927 249
989 249
989 286
979 286
1 0 12 0 0 4096 0 6 0 0 23 4
980 230
993 230
993 231
998 231
2 2 13 0 0 12416 0 7 43 0 0 6
653 215
641 215
641 241
703 241
703 276
687 276
1 0 14 0 0 4096 0 7 0 0 24 2
689 215
712 215
2 2 15 0 0 12416 0 8 38 0 0 6
372 220
361 220
361 240
419 240
419 275
414 275
1 0 16 0 0 4096 0 8 0 0 25 2
408 220
425 220
2 2 17 0 0 12416 0 9 33 0 0 6
126 217
111 217
111 236
173 236
173 265
156 265
1 0 18 0 0 4096 0 9 0 0 26 2
162 217
183 217
1 2 12 0 0 4224 0 19 26 0 0 4
998 179
998 254
1064 254
1064 263
1 2 14 0 0 4224 0 21 45 0 0 4
712 179
712 246
765 246
765 259
1 2 16 0 0 4224 0 23 36 0 0 4
425 176
425 242
485 242
485 255
1 2 18 0 0 4224 0 25 31 0 0 4
183 177
183 240
235 240
235 253
1 0 19 0 0 4096 0 1 0 0 55 3
1165 346
1165 337
1081 337
2 0 2 0 0 0 0 10 0 0 31 4
43 485
43 541
259 541
259 515
3 1 20 0 0 8320 0 35 10 0 0 3
46 323
43 323
43 465
2 0 2 0 0 0 0 13 0 0 31 2
508 478
508 515
2 1 2 0 0 0 0 12 11 0 0 4
258 490
258 515
629 515
629 573
3 1 21 0 0 4224 0 27 15 0 0 4
1074 404
1074 476
1076 476
1076 484
3 1 22 0 0 4224 0 44 14 0 0 2
788 396
788 463
3 1 23 0 0 4224 0 37 13 0 0 2
508 392
508 458
3 1 24 0 0 4224 0 32 12 0 0 2
258 390
258 470
3 0 2 0 0 0 0 25 0 0 43 2
179 143
179 122
3 0 2 0 0 0 0 24 0 0 43 2
269 146
269 122
3 0 2 0 0 0 0 23 0 0 43 2
421 142
421 122
3 0 2 0 0 0 0 22 0 0 43 2
519 142
519 122
3 0 2 0 0 0 0 21 0 0 43 2
708 145
708 122
3 0 2 0 0 0 0 20 0 0 43 2
791 146
791 122
3 0 2 0 0 0 0 19 0 0 43 2
994 145
994 122
1 3 2 0 0 8320 0 16 18 0 0 4
78 126
78 122
1085 122
1085 144
2 0 25 0 0 4096 9 25 0 0 51 2
187 143
187 100
2 0 25 0 0 0 9 24 0 0 51 4
277 146
277 134
278 134
278 100
2 0 25 0 0 0 9 23 0 0 51 2
429 142
429 100
2 0 25 0 0 0 9 22 0 0 51 2
527 142
527 100
2 0 25 0 0 4096 9 21 0 0 51 2
716 145
716 100
2 0 25 0 0 4096 9 20 0 0 51 2
799 146
799 100
2 0 25 0 0 0 9 19 0 0 51 4
1002 145
1002 134
1003 134
1003 100
1 2 25 0 0 8320 9 17 18 0 0 4
120 71
120 100
1093 100
1093 144
3 0 26 0 0 4096 0 40 0 0 60 2
296 325
267 325
3 0 27 0 0 4096 0 41 0 0 65 2
576 329
517 329
3 0 28 0 0 4096 0 30 0 0 66 2
862 337
797 337
1 1 19 0 0 8320 0 29 27 0 0 5
983 427
1032 427
1032 337
1083 337
1083 355
3 1 29 0 0 8320 0 29 30 0 0 4
938 418
930 418
930 346
908 346
3 2 30 0 0 8320 0 28 30 0 0 4
934 295
930 295
930 328
908 328
1 0 31 0 0 8192 16 28 0 0 59 4
979 304
1035 304
1035 240
1089 240
1 1 31 0 0 4224 16 18 26 0 0 4
1089 178
1089 254
1082 254
1082 263
1 1 26 0 0 8320 0 34 32 0 0 5
182 420
213 420
213 307
267 307
267 341
3 1 32 0 0 8320 0 34 35 0 0 4
137 411
114 411
114 332
92 332
3 2 33 0 0 8320 0 33 35 0 0 4
111 274
102 274
102 314
92 314
1 0 34 0 0 12416 21 33 0 0 64 4
156 283
212 283
212 226
273 226
1 1 34 0 0 0 21 24 31 0 0 4
273 180
273 240
253 240
253 253
1 1 27 0 0 8320 0 39 37 0 0 5
421 411
466 411
466 325
517 325
517 343
1 1 28 0 0 8320 0 42 44 0 0 5
707 414
743 414
743 313
797 313
797 347
3 1 35 0 0 8320 0 39 40 0 0 4
376 402
364 402
364 334
342 334
3 2 36 0 0 8320 0 38 40 0 0 4
369 284
364 284
364 316
342 316
1 0 37 0 0 8192 26 38 0 0 70 4
414 293
467 293
467 228
523 228
1 1 37 0 0 4224 26 22 36 0 0 4
523 176
523 242
503 242
503 255
3 1 38 0 0 8320 0 42 41 0 0 4
662 405
644 405
644 338
622 338
3 2 39 0 0 8320 0 43 41 0 0 4
642 285
633 285
633 320
622 320
1 0 40 0 0 8192 30 43 0 0 74 4
687 294
748 294
748 232
795 232
1 1 40 0 0 4224 30 20 45 0 0 4
795 180
795 246
783 246
783 259
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
