CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
10 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
58 C:\Users\joaop\Desktop\circuitmaker+traxmaker+2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
41
2 +V
167 1174 334 0 1 3
0 0
0
0 0 54240 0
3 10V
-11 -22 10 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
828 0 0
2
42691.7 0
0
9 Inverter~
13 1004 223 0 1 22
0 0
0
0 0 608 270
6 74LS04
-21 -19 21 -11
3 U6D
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 6 0
1 U
6187 0 0
2
42691.7 0
0
9 Inverter~
13 718 219 0 1 22
0 0
0
0 0 608 270
6 74LS04
-21 -19 21 -11
3 U6C
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 6 0
1 U
7107 0 0
2
42691.7 0
0
9 Inverter~
13 431 215 0 1 22
0 0
0
0 0 608 270
6 74LS04
-21 -19 21 -11
3 U6B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 6 0
1 U
6433 0 0
2
42691.7 0
0
9 Inverter~
13 189 212 0 1 22
0 0
0
0 0 608 270
6 74LS04
-21 -19 21 -11
3 U6A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 6 0
1 U
8559 0 0
2
42691.7 0
0
6 74136~
219 780 284 0 3 22
0 22 22 29
0
0 0 608 270
7 74LS136
-24 -24 25 -16
3 U4D
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
3674 0 0
2
42691.7 36
0
6 74136~
219 794 372 0 3 22
0 12 29 6
0
0 0 608 270
7 74LS136
-24 -24 25 -16
3 U4C
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
5697 0 0
2
42691.7 35
0
9 2-In AND~
219 684 284 0 3 22
0 22 22 28
0
0 0 608 180
6 74LS08
-21 -24 21 -16
3 U5D
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
3805 0 0
2
42691.7 33
0
9 2-In AND~
219 700 381 0 3 22
0 12 29 27
0
0 0 608 180
6 74LS08
-21 -24 21 -16
3 U5C
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
5219 0 0
2
42691.7 32
0
8 2-In OR~
219 612 335 0 3 22
0 27 28 11
0
0 0 608 180
6 74LS32
-21 -24 21 -16
3 U3D
1 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
3795 0 0
2
42691.7 31
0
8 2-In OR~
219 332 331 0 3 22
0 23 24 10
0
0 0 608 180
6 74LS32
-21 -24 21 -16
3 U3C
1 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
3637 0 0
2
42691.7 30
0
9 2-In AND~
219 420 377 0 3 22
0 11 25 23
0
0 0 608 180
6 74LS08
-21 -24 21 -16
3 U5B
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
3226 0 0
2
42691.7 29
0
9 2-In AND~
219 404 280 0 3 22
0 22 22 24
0
0 0 608 180
6 74LS08
-21 -24 21 -16
3 U5A
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
6966 0 0
2
42691.7 28
0
6 74136~
219 514 368 0 3 22
0 11 25 7
0
0 0 608 270
7 74LS136
-24 -24 25 -16
3 U4B
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
9796 0 0
2
42691.7 27
0
6 74136~
219 500 280 0 3 22
0 22 22 25
0
0 0 608 270
7 74LS136
-24 -24 25 -16
3 U4A
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
5952 0 0
2
42691.7 26
0
8 2-In OR~
219 82 329 0 3 22
0 18 19 4
0
0 0 608 180
6 74LS32
-21 -24 21 -16
3 U3B
1 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
3649 0 0
2
42691.7 25
0
9 2-In AND~
219 170 375 0 3 22
0 10 20 18
0
0 0 608 180
6 74LS08
-21 -24 21 -16
3 U2D
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
3716 0 0
2
42691.7 24
0
9 2-In AND~
219 154 278 0 3 22
0 22 22 19
0
0 0 608 180
6 74LS08
-21 -24 21 -16
3 U2C
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
4797 0 0
2
42691.7 23
0
6 74136~
219 264 366 0 3 22
0 10 20 8
0
0 0 608 270
7 74LS136
-24 -24 25 -16
3 U1D
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
4681 0 0
2
42691.7 22
0
6 74136~
219 250 278 0 3 22
0 22 22 20
0
0 0 608 270
7 74LS136
-24 -24 25 -16
3 U1C
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
9730 0 0
2
42691.7 21
0
8 2-In OR~
219 898 343 0 3 22
0 13 14 12
0
0 0 608 180
6 74LS32
-21 -24 21 -16
3 U3A
1 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
9874 0 0
2
42691.7 20
0
9 2-In AND~
219 986 389 0 3 22
0 2 15 13
0
0 0 608 180
6 74LS08
-21 -24 21 -16
3 U2B
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
364 0 0
2
42691.7 19
0
9 2-In AND~
219 970 292 0 3 22
0 22 22 14
0
0 0 608 180
6 74LS08
-21 -24 21 -16
3 U2A
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3656 0 0
2
42691.7 18
0
6 74136~
219 1080 380 0 3 22
0 2 15 5
0
0 0 608 270
7 74LS136
-24 -24 25 -16
3 U1B
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
3131 0 0
2
42691.7 17
0
6 74136~
219 1066 292 0 3 22
0 22 22 15
0
0 0 608 270
7 74LS136
-24 -24 25 -16
3 U1A
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
6772 0 0
2
42691.7 16
0
12 SPDT Switch~
164 193 165 0 10 11
0 22 22 2 0 0 0 0 0 0
1
0
0 0 4704 270
0
2 S1
9 -4 23 4
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
9557 0 0
2
42691.7 15
0
12 SPDT Switch~
164 283 168 0 10 11
0 22 22 2 0 0 0 0 0 0
1
0
0 0 4704 270
0
2 S2
9 -4 23 4
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
5789 0 0
2
42691.7 14
0
12 SPDT Switch~
164 435 164 0 10 11
0 22 22 2 0 0 0 0 0 0
1
0
0 0 4704 270
0
2 S3
9 -4 23 4
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
7328 0 0
2
42691.7 13
0
12 SPDT Switch~
164 533 164 0 10 11
0 22 22 2 0 0 0 0 0 0
1
0
0 0 4704 270
0
2 S4
9 -4 23 4
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
4799 0 0
2
42691.7 12
0
12 SPDT Switch~
164 722 167 0 10 11
0 22 22 2 0 0 0 0 0 0
1
0
0 0 4704 270
0
2 S5
9 -4 23 4
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
9196 0 0
2
42691.7 11
0
12 SPDT Switch~
164 805 168 0 10 11
0 22 22 2 0 0 0 0 0 0
1
0
0 0 4704 270
0
2 S6
9 -4 23 4
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
3857 0 0
2
42691.7 10
0
12 SPDT Switch~
164 1008 167 0 10 11
0 22 22 2 0 0 0 0 0 0
1
0
0 0 4704 270
0
2 S7
9 -4 23 4
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
7125 0 0
2
42691.7 9
0
12 SPDT Switch~
164 1099 166 0 10 11
0 22 22 2 0 0 0 0 0 0
1
0
0 0 4704 270
0
2 S8
9 -4 23 4
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
3641 0 0
2
42691.7 8
0
2 +V
167 129 68 0 1 3
0 22
0
0 0 54240 0
3 10V
-11 -23 10 -15
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9821 0 0
2
42691.7 7
0
7 Ground~
168 87 138 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3187 0 0
2
42691.7 6
0
4 LED~
171 1085 500 0 1 2
10 5
0
0 0 880 0
4 LED0
17 0 45 8
2 D1
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
762 0 0
2
42691.7 5
0
4 LED~
171 804 491 0 1 2
10 6
0
0 0 880 0
4 LED0
17 0 45 8
2 D2
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
39 0 0
2
42691.7 4
0
4 LED~
171 517 474 0 1 2
10 7
0
0 0 880 0
4 LED0
17 0 45 8
2 D3
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
9450 0 0
2
42691.7 3
0
4 LED~
171 267 486 0 1 2
10 8
0
0 0 880 0
4 LED0
17 0 45 8
2 D4
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3236 0 0
2
42691.7 2
0
7 Ground~
168 638 585 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3321 0 0
2
42691.7 1
0
4 LED~
171 52 481 0 1 2
10 4
0
0 0 880 0
4 LED0
17 0 45 8
2 D5
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
8879 0 0
2
42691.7 0
0
70
1 0 0 0 0 0 0 1 0 0 43 2
1174 343
1090 343
2 0 0 0 0 0 0 23 0 0 9 4
988 283
1002 283
1002 257
1007 257
2 0 0 0 0 0 0 8 0 0 8 4
702 275
716 275
716 252
721 252
2 0 0 0 0 0 0 13 0 0 7 4
422 271
429 271
429 247
434 247
2 0 0 0 0 0 0 18 0 0 6 4
172 269
187 269
187 245
192 245
2 2 0 0 0 0 0 5 20 0 0 4
192 230
192 246
244 246
244 259
2 2 0 0 0 0 0 4 15 0 0 4
434 233
434 248
494 248
494 261
2 2 0 0 0 0 0 3 6 0 0 4
721 237
721 252
774 252
774 265
2 2 0 0 0 0 0 2 25 0 0 4
1007 241
1007 260
1060 260
1060 273
1 1 0 0 0 0 0 26 5 0 0 2
192 183
192 194
1 1 0 0 0 0 0 32 2 0 0 2
1007 185
1007 205
1 1 0 0 0 0 0 30 3 0 0 2
721 185
721 201
1 1 0 0 0 0 0 28 4 0 0 2
434 182
434 197
2 0 2 0 0 0 0 41 0 0 19 3
52 491
52 544
277 544
3 1 4 0 0 0 0 16 41 0 0 3
55 329
52 329
52 471
2 0 2 0 0 0 0 38 0 0 19 2
517 484
517 544
2 0 2 0 0 0 0 37 0 0 18 2
804 501
804 544
2 1 2 0 0 0 0 36 40 0 0 4
1085 510
1085 544
638 544
638 579
2 1 2 0 0 0 0 39 40 0 0 4
267 496
267 544
638 544
638 579
3 1 5 0 0 0 0 24 36 0 0 4
1083 410
1083 482
1085 482
1085 490
3 1 6 0 0 0 0 7 37 0 0 4
797 402
797 473
804 473
804 481
3 1 7 0 0 0 0 14 38 0 0 2
517 398
517 464
3 1 8 0 0 0 0 19 39 0 0 2
267 396
267 476
3 0 2 0 0 0 0 26 0 0 31 2
188 149
188 128
3 0 2 0 0 0 0 27 0 0 31 2
278 152
278 128
3 0 2 0 0 0 0 28 0 0 31 2
430 148
430 128
3 0 2 0 0 0 0 29 0 0 31 2
528 148
528 128
3 0 2 0 0 0 0 30 0 0 31 2
717 151
717 128
3 0 2 0 0 0 0 31 0 0 31 2
800 152
800 128
3 0 2 0 0 0 0 32 0 0 31 2
1003 151
1003 128
1 3 2 0 0 0 0 35 33 0 0 4
87 132
87 128
1094 128
1094 150
2 0 22 0 0 0 9 26 0 0 39 2
196 149
196 106
2 0 22 0 0 0 9 27 0 0 39 4
286 152
286 140
287 140
287 106
2 0 22 0 0 0 9 28 0 0 39 2
438 148
438 106
2 0 22 0 0 0 9 29 0 0 39 2
536 148
536 106
2 0 22 0 0 0 9 30 0 0 39 2
725 151
725 106
2 0 22 0 0 0 9 31 0 0 39 2
808 152
808 106
2 0 22 0 0 0 9 32 0 0 39 4
1011 151
1011 140
1012 140
1012 106
1 2 22 0 0 0 9 34 33 0 0 4
129 77
129 106
1102 106
1102 150
3 0 10 0 0 0 0 11 0 0 50 2
305 331
276 331
3 0 11 0 0 0 0 10 0 0 57 2
585 335
526 335
3 0 12 0 0 0 0 21 0 0 58 2
871 343
806 343
1 1 2 0 0 0 0 22 24 0 0 5
1004 398
1041 398
1041 343
1092 343
1092 361
3 1 13 0 0 0 0 22 21 0 0 4
959 389
939 389
939 352
917 352
3 2 14 0 0 0 0 23 21 0 0 4
943 292
939 292
939 334
917 334
3 0 15 0 0 0 0 25 0 0 47 3
1069 322
1069 348
1055 348
2 2 15 0 0 0 0 22 24 0 0 5
1004 380
1055 380
1055 348
1074 348
1074 361
1 0 22 0 0 0 16 23 0 0 49 4
988 301
1044 301
1044 246
1098 246
1 1 22 0 0 0 16 33 25 0 0 4
1098 184
1098 260
1078 260
1078 273
1 1 10 0 0 0 0 17 19 0 0 5
188 384
225 384
225 329
276 329
276 347
3 1 18 0 0 0 0 17 16 0 0 4
143 375
123 375
123 338
101 338
3 2 19 0 0 0 0 18 16 0 0 4
127 278
123 278
123 320
101 320
3 0 20 0 0 16 0 20 0 0 54 3
253 308
245 308
245 340
2 2 20 0 0 0 0 17 19 0 0 5
188 366
245 366
245 340
258 340
258 347
1 0 22 0 0 0 21 18 0 0 56 4
172 287
221 287
221 232
282 232
1 1 22 0 0 0 21 27 20 0 0 4
282 186
282 246
262 246
262 259
1 1 11 0 0 0 0 12 14 0 0 5
438 386
475 386
475 331
526 331
526 349
1 1 12 0 0 0 0 9 7 0 0 5
718 390
749 390
749 335
806 335
806 353
3 1 23 0 0 0 0 12 11 0 0 4
393 377
373 377
373 340
351 340
3 2 24 0 0 0 0 13 11 0 0 4
377 280
373 280
373 322
351 322
3 0 25 0 0 0 0 15 0 0 62 3
503 310
503 336
488 336
2 2 25 0 0 0 0 12 14 0 0 5
438 368
488 368
488 336
508 336
508 349
1 0 22 0 0 0 26 13 0 0 64 4
422 289
476 289
476 234
532 234
1 1 22 0 0 0 26 29 15 0 0 4
532 182
532 248
512 248
512 261
3 1 27 0 0 0 0 9 10 0 0 4
673 381
653 381
653 344
631 344
3 2 28 0 0 0 0 8 10 0 0 4
657 284
653 284
653 326
631 326
3 0 29 0 0 0 0 6 0 0 68 3
783 314
783 340
765 340
2 2 29 0 0 0 0 9 7 0 0 5
718 372
765 372
765 340
788 340
788 353
1 0 22 0 0 0 30 8 0 0 70 4
702 293
757 293
757 238
804 238
1 1 22 0 0 0 30 31 6 0 0 4
804 186
804 252
792 252
792 265
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
