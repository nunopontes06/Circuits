CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
130 40 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
58 C:\Users\joaop\Desktop\circuitmaker+traxmaker+2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
37
4 LED~
171 152 474 0 2 2
10 4 2
0
0 0 864 0
4 LED0
17 0 45 8
2 D5
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
9968 0 0
2
5.89777e-315 0
0
7 Ground~
168 738 578 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9281 0 0
2
5.89777e-315 0
0
4 LED~
171 377 479 0 2 2
10 8 2
0
0 0 864 0
4 LED0
17 0 45 8
2 D4
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
8464 0 0
2
5.89777e-315 0
0
4 LED~
171 617 467 0 2 2
10 7 2
0
0 0 864 0
4 LED0
17 0 45 8
2 D3
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
7168 0 0
2
5.89777e-315 0
0
4 LED~
171 904 484 0 2 2
10 6 2
0
0 0 864 0
4 LED0
17 0 45 8
2 D2
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3171 0 0
2
5.89777e-315 0
0
4 LED~
171 1185 493 0 2 2
10 5 2
0
0 0 864 0
4 LED0
17 0 45 8
2 D1
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
4139 0 0
2
5.89777e-315 0
0
7 Ground~
168 187 131 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6435 0 0
2
5.89777e-315 0
0
2 +V
167 229 61 0 1 3
0 22
0
0 0 54256 0
3 10V
-11 -23 10 -15
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5283 0 0
2
5.89777e-315 0
0
12 SPDT Switch~
164 1199 159 0 10 11
0 22 22 2 0 0 0 0 0 0
1
0
0 0 4720 270
0
2 S8
9 -4 23 4
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
6874 0 0
2
5.89777e-315 0
0
12 SPDT Switch~
164 1108 160 0 10 11
0 22 22 2 0 0 0 0 0 0
1
0
0 0 4720 270
0
2 S7
9 -4 23 4
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
5305 0 0
2
5.89777e-315 0
0
12 SPDT Switch~
164 905 161 0 10 11
0 22 22 2 0 0 0 0 0 0
1
0
0 0 4720 270
0
2 S6
9 -4 23 4
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
34 0 0
2
5.89777e-315 0
0
12 SPDT Switch~
164 822 160 0 10 11
0 22 22 2 0 0 0 0 0 0
1
0
0 0 4720 270
0
2 S5
9 -4 23 4
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
969 0 0
2
5.89777e-315 0
0
12 SPDT Switch~
164 633 157 0 10 11
0 22 22 2 0 0 0 0 0 0
1
0
0 0 4720 270
0
2 S4
9 -4 23 4
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
8402 0 0
2
5.89777e-315 0
0
12 SPDT Switch~
164 535 157 0 10 11
0 22 22 2 0 0 0 0 0 0
1
0
0 0 4720 270
0
2 S3
9 -4 23 4
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
3751 0 0
2
5.89777e-315 0
0
12 SPDT Switch~
164 383 161 0 10 11
0 22 22 2 0 0 0 0 0 0
1
0
0 0 4720 270
0
2 S2
9 -4 23 4
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
4292 0 0
2
5.89777e-315 0
0
12 SPDT Switch~
164 293 158 0 10 11
0 22 22 2 0 0 0 0 0 0
1
0
0 0 4720 270
0
2 S1
9 -4 23 4
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
6118 0 0
2
5.89777e-315 0
0
6 74136~
219 1166 285 0 3 22
0 22 22 15
0
0 0 624 270
7 74LS136
-24 -24 25 -16
3 U5D
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
34 0 0
2
5.89777e-315 5.34643e-315
0
6 74136~
219 1180 373 0 3 22
0 2 15 5
0
0 0 624 270
7 74LS136
-24 -24 25 -16
3 U5C
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
6357 0 0
2
5.89777e-315 5.32571e-315
0
9 2-In AND~
219 1070 285 0 3 22
0 22 22 14
0
0 0 624 180
6 74LS08
-21 -24 21 -16
3 U4D
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
319 0 0
2
5.89777e-315 5.30499e-315
0
9 2-In AND~
219 1086 382 0 3 22
0 2 15 13
0
0 0 624 180
6 74LS08
-21 -24 21 -16
3 U4C
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
3976 0 0
2
5.89777e-315 5.26354e-315
0
8 2-In OR~
219 998 336 0 3 22
0 13 14 12
0
0 0 624 180
6 74LS32
-21 -24 21 -16
3 U3D
1 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
7634 0 0
2
5.89777e-315 0
0
6 74136~
219 350 271 0 3 22
0 22 22 20
0
0 0 624 270
7 74LS136
-24 -24 25 -16
3 U5B
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
523 0 0
2
5.89777e-315 5.34643e-315
0
6 74136~
219 364 359 0 3 22
0 10 20 8
0
0 0 624 270
7 74LS136
-24 -24 25 -16
3 U5A
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
6748 0 0
2
5.89777e-315 5.32571e-315
0
9 2-In AND~
219 254 271 0 3 22
0 22 22 19
0
0 0 624 180
6 74LS08
-21 -24 21 -16
3 U4B
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
6901 0 0
2
5.89777e-315 5.30499e-315
0
9 2-In AND~
219 270 368 0 3 22
0 10 20 18
0
0 0 624 180
6 74LS08
-21 -24 21 -16
3 U4A
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
842 0 0
2
5.89777e-315 5.26354e-315
0
8 2-In OR~
219 182 322 0 3 22
0 18 19 4
0
0 0 624 180
6 74LS32
-21 -24 21 -16
3 U3C
1 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
3277 0 0
2
5.89777e-315 0
0
6 74136~
219 600 273 0 3 22
0 22 22 25
0
0 0 624 270
7 74LS136
-24 -24 25 -16
3 U1D
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
4212 0 0
2
5.89777e-315 5.34643e-315
0
6 74136~
219 614 361 0 3 22
0 11 25 7
0
0 0 624 270
7 74LS136
-24 -24 25 -16
3 U1C
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
4720 0 0
2
5.89777e-315 5.32571e-315
0
9 2-In AND~
219 504 273 0 3 22
0 22 22 24
0
0 0 624 180
6 74LS08
-21 -24 21 -16
3 U2D
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
5551 0 0
2
5.89777e-315 5.30499e-315
0
9 2-In AND~
219 520 370 0 3 22
0 11 25 23
0
0 0 624 180
6 74LS08
-21 -24 21 -16
3 U2C
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
6986 0 0
2
5.89777e-315 5.26354e-315
0
8 2-In OR~
219 432 324 0 3 22
0 23 24 10
0
0 0 624 180
6 74LS32
-21 -24 21 -16
3 U3B
1 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
8745 0 0
2
5.89777e-315 0
0
8 2-In OR~
219 712 328 0 3 22
0 27 28 11
0
0 0 624 180
6 74LS32
-21 -24 21 -16
3 U3A
1 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
9592 0 0
2
5.89777e-315 0
0
9 2-In AND~
219 800 374 0 3 22
0 12 29 27
0
0 0 624 180
6 74LS08
-21 -24 21 -16
3 U2B
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
8748 0 0
2
5.89777e-315 0
0
9 2-In AND~
219 784 277 0 3 22
0 22 22 28
0
0 0 624 180
6 74LS08
-21 -24 21 -16
3 U2A
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
7168 0 0
2
5.89777e-315 0
0
7 Ground~
168 1311 363 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
631 0 0
2
5.89777e-315 0
0
6 74136~
219 894 365 0 3 22
0 12 29 6
0
0 0 624 270
7 74LS136
-24 -24 25 -16
3 U1B
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
9466 0 0
2
5.89777e-315 0
0
6 74136~
219 880 277 0 3 22
0 22 22 29
0
0 0 624 270
7 74LS136
-24 -24 25 -16
3 U1A
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3266 0 0
2
5.89777e-315 0
0
66
2 0 22 0 0 8192 3 29 0 0 2 4
522 264
529 264
529 241
534 241
1 2 22 0 0 4224 3 14 27 0 0 4
534 175
534 241
594 241
594 254
2 0 2 0 0 8192 0 1 0 0 8 3
152 484
152 537
377 537
3 1 4 0 0 8320 0 26 1 0 0 3
155 322
152 322
152 464
2 0 2 0 0 0 0 4 0 0 8 2
617 477
617 537
2 0 2 0 0 0 0 5 0 0 7 2
904 494
904 537
2 1 2 0 0 8192 0 6 2 0 0 4
1185 503
1185 537
738 537
738 572
2 1 2 0 0 0 0 3 2 0 0 4
377 489
377 537
738 537
738 572
3 1 5 0 0 4224 0 18 6 0 0 4
1183 403
1183 475
1185 475
1185 483
3 1 6 0 0 4224 0 36 5 0 0 4
897 395
897 466
904 466
904 474
3 1 7 0 0 4224 0 28 4 0 0 2
617 391
617 457
3 1 8 0 0 4224 0 23 3 0 0 4
367 389
367 461
377 461
377 469
3 0 2 0 0 0 0 16 0 0 20 2
288 142
288 121
3 0 2 0 0 0 0 15 0 0 20 2
378 145
378 121
3 0 2 0 0 0 0 14 0 0 20 2
530 141
530 121
3 0 2 0 0 0 0 13 0 0 20 2
628 141
628 121
3 0 2 0 0 0 0 12 0 0 20 2
817 144
817 121
3 0 2 0 0 0 0 11 0 0 20 2
900 145
900 121
3 0 2 0 0 0 0 10 0 0 20 2
1103 144
1103 121
1 3 2 0 0 8320 0 7 9 0 0 4
187 125
187 121
1194 121
1194 143
2 0 22 0 0 4096 9 16 0 0 28 2
296 142
296 99
2 0 22 0 0 0 9 15 0 0 28 4
386 145
386 133
387 133
387 99
2 0 22 0 0 0 9 14 0 0 28 2
538 141
538 99
2 0 22 0 0 0 9 13 0 0 28 2
636 141
636 99
2 0 22 0 0 4096 9 12 0 0 28 2
825 144
825 99
2 0 22 0 0 4096 9 11 0 0 28 2
908 145
908 99
2 0 22 0 0 0 9 10 0 0 28 4
1111 144
1111 133
1112 133
1112 99
1 2 22 0 0 8320 9 8 9 0 0 4
229 70
229 99
1202 99
1202 143
1 0 2 0 0 0 0 35 0 0 33 3
1311 357
1311 344
1192 344
3 0 10 0 0 4096 0 31 0 0 42 2
405 324
376 324
3 0 11 0 0 4224 0 32 0 0 51 2
685 328
626 328
3 0 12 0 0 4224 0 21 0 0 52 2
971 336
906 336
1 1 2 0 0 0 0 20 18 0 0 5
1104 391
1141 391
1141 336
1192 336
1192 354
3 1 13 0 0 8320 0 20 21 0 0 4
1059 382
1039 382
1039 345
1017 345
3 2 14 0 0 8320 0 19 21 0 0 4
1043 285
1039 285
1039 327
1017 327
3 0 15 0 0 4096 0 17 0 0 37 3
1169 315
1169 341
1155 341
2 2 15 0 0 4224 0 20 18 0 0 5
1104 373
1155 373
1155 341
1174 341
1174 354
1 0 22 0 0 4096 16 19 0 0 40 4
1088 294
1144 294
1144 239
1198 239
2 0 22 0 0 8192 17 19 0 0 41 4
1088 276
1103 276
1103 244
1107 244
1 1 22 0 0 4224 16 9 17 0 0 4
1198 177
1198 253
1178 253
1178 266
1 2 22 0 0 4224 17 10 17 0 0 4
1107 178
1107 253
1160 253
1160 266
1 1 10 0 0 8320 0 25 23 0 0 5
288 377
328 377
328 322
376 322
376 340
3 1 18 0 0 8320 0 25 26 0 0 4
243 368
223 368
223 331
201 331
3 2 19 0 0 8320 0 24 26 0 0 4
227 271
223 271
223 313
201 313
3 0 20 0 0 4096 0 22 0 0 46 3
353 301
353 327
340 327
2 2 20 0 0 4224 0 25 23 0 0 5
288 359
340 359
340 327
358 327
358 340
1 0 22 0 0 12416 21 24 0 0 49 4
272 280
321 280
321 225
382 225
2 0 22 0 0 8192 0 24 0 0 50 4
272 262
287 262
287 230
292 230
1 1 22 0 0 0 21 15 22 0 0 4
382 179
382 239
362 239
362 252
1 2 22 0 0 4224 0 16 22 0 0 4
292 176
292 239
344 239
344 252
1 1 11 0 0 128 0 30 28 0 0 5
538 379
575 379
575 324
626 324
626 342
1 1 12 0 0 16 0 33 36 0 0 5
818 383
849 383
849 328
906 328
906 346
3 1 23 0 0 8320 0 30 31 0 0 4
493 370
473 370
473 333
451 333
3 2 24 0 0 8320 0 29 31 0 0 4
477 273
473 273
473 315
451 315
3 0 25 0 0 4096 0 27 0 0 56 3
603 303
603 329
588 329
2 2 25 0 0 4224 0 30 28 0 0 5
538 361
588 361
588 329
608 329
608 342
1 0 22 0 0 12416 26 29 0 0 58 4
522 282
576 282
576 227
632 227
1 1 22 0 0 4224 26 13 27 0 0 4
632 175
632 241
612 241
612 254
3 1 27 0 0 8320 0 33 32 0 0 4
773 374
753 374
753 337
731 337
3 2 28 0 0 8320 0 34 32 0 0 4
757 277
753 277
753 319
731 319
3 0 29 0 0 4096 0 37 0 0 62 3
883 307
883 333
865 333
2 2 29 0 0 4224 0 33 36 0 0 5
818 365
865 365
865 333
888 333
888 346
1 0 22 0 0 4224 30 34 0 0 65 4
802 286
857 286
857 231
904 231
2 0 22 0 0 8192 31 34 0 0 66 4
802 268
817 268
817 236
821 236
1 1 22 0 0 4224 30 11 37 0 0 4
904 179
904 245
892 245
892 258
1 2 22 0 0 4224 31 12 37 0 0 4
821 178
821 245
874 245
874 258
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
